library ieee;
use ieee.std_logic_1164.all;

entity wave_lut is
    generic (
        signal_width: integer := 8
    );
    port (
		index : in std_logic_vector(15 downto 0);
		output : out std_logic_vector(signal_width - 1 downto 0)
    );
end;

architecture behavior of wave_lut is

begin

process (index)
begin

case index(9 downto 0) is

-- sine wave
when "0000000000" => output <= "00000000";
when "0000000001" => output <= "00000011";
when "0000000010" => output <= "00000110";
when "0000000011" => output <= "00001001";
when "0000000100" => output <= "00001100";
when "0000000101" => output <= "00001111";
when "0000000110" => output <= "00010010";
when "0000000111" => output <= "00010101";
when "0000001000" => output <= "00011001";
when "0000001001" => output <= "00011100";
when "0000001010" => output <= "00011111";
when "0000001011" => output <= "00100010";
when "0000001100" => output <= "00100101";
when "0000001101" => output <= "00101000";
when "0000001110" => output <= "00101011";
when "0000001111" => output <= "00101110";
when "0000010000" => output <= "00110001";
when "0000010001" => output <= "00110100";
when "0000010010" => output <= "00110110";
when "0000010011" => output <= "00111001";
when "0000010100" => output <= "00111100";
when "0000010101" => output <= "00111111";
when "0000010110" => output <= "01000010";
when "0000010111" => output <= "01000100";
when "0000011000" => output <= "01000111";
when "0000011001" => output <= "01001001";
when "0000011010" => output <= "01001100";
when "0000011011" => output <= "01001111";
when "0000011100" => output <= "01010001";
when "0000011101" => output <= "01010011";
when "0000011110" => output <= "01010110";
when "0000011111" => output <= "01011000";
when "0000100000" => output <= "01011010";
when "0000100001" => output <= "01011100";
when "0000100010" => output <= "01011111";
when "0000100011" => output <= "01100001";
when "0000100100" => output <= "01100011";
when "0000100101" => output <= "01100101";
when "0000100110" => output <= "01100111";
when "0000100111" => output <= "01101000";
when "0000101000" => output <= "01101010";
when "0000101001" => output <= "01101100";
when "0000101010" => output <= "01101110";
when "0000101011" => output <= "01101111";
when "0000101100" => output <= "01110001";
when "0000101101" => output <= "01110010";
when "0000101110" => output <= "01110011";
when "0000101111" => output <= "01110101";
when "0000110000" => output <= "01110110";
when "0000110001" => output <= "01110111";
when "0000110010" => output <= "01111000";
when "0000110011" => output <= "01111001";
when "0000110100" => output <= "01111010";
when "0000110101" => output <= "01111011";
when "0000110110" => output <= "01111100";
when "0000110111" => output <= "01111101";
when "0000111000" => output <= "01111101";
when "0000111001" => output <= "01111110";
when "0000111010" => output <= "01111110";
when "0000111011" => output <= "01111111";
when "0000111100" => output <= "01111111";
when "0000111101" => output <= "01111111";
when "0000111110" => output <= "01111111";
when "0000111111" => output <= "01111111";
when "0001000000" => output <= "01111111";
when "0001000001" => output <= "01111111";
when "0001000010" => output <= "01111111";
when "0001000011" => output <= "01111111";
when "0001000100" => output <= "01111111";
when "0001000101" => output <= "01111110";
when "0001000110" => output <= "01111110";
when "0001000111" => output <= "01111101";
when "0001001000" => output <= "01111101";
when "0001001001" => output <= "01111100";
when "0001001010" => output <= "01111011";
when "0001001011" => output <= "01111011";
when "0001001100" => output <= "01111010";
when "0001001101" => output <= "01111001";
when "0001001110" => output <= "01111000";
when "0001001111" => output <= "01110111";
when "0001010000" => output <= "01110101";
when "0001010001" => output <= "01110100";
when "0001010010" => output <= "01110011";
when "0001010011" => output <= "01110001";
when "0001010100" => output <= "01110000";
when "0001010101" => output <= "01101110";
when "0001010110" => output <= "01101101";
when "0001010111" => output <= "01101011";
when "0001011000" => output <= "01101001";
when "0001011001" => output <= "01101000";
when "0001011010" => output <= "01100110";
when "0001011011" => output <= "01100100";
when "0001011100" => output <= "01100010";
when "0001011101" => output <= "01100000";
when "0001011110" => output <= "01011110";
when "0001011111" => output <= "01011011";
when "0001100000" => output <= "01011001";
when "0001100001" => output <= "01010111";
when "0001100010" => output <= "01010101";
when "0001100011" => output <= "01010010";
when "0001100100" => output <= "01010000";
when "0001100101" => output <= "01001101";
when "0001100110" => output <= "01001011";
when "0001100111" => output <= "01001000";
when "0001101000" => output <= "01000110";
when "0001101001" => output <= "01000011";
when "0001101010" => output <= "01000000";
when "0001101011" => output <= "00111101";
when "0001101100" => output <= "00111011";
when "0001101101" => output <= "00111000";
when "0001101110" => output <= "00110101";
when "0001101111" => output <= "00110010";
when "0001110000" => output <= "00101111";
when "0001110001" => output <= "00101100";
when "0001110010" => output <= "00101001";
when "0001110011" => output <= "00100110";
when "0001110100" => output <= "00100011";
when "0001110101" => output <= "00100000";
when "0001110110" => output <= "00011101";
when "0001110111" => output <= "00011010";
when "0001111000" => output <= "00010111";
when "0001111001" => output <= "00010100";
when "0001111010" => output <= "00010001";
when "0001111011" => output <= "00001110";
when "0001111100" => output <= "00001011";
when "0001111101" => output <= "00000111";
when "0001111110" => output <= "00000100";
when "0001111111" => output <= "00000001";
when "0010000000" => output <= "11111111";
when "0010000001" => output <= "11111100";
when "0010000010" => output <= "11111001";
when "0010000011" => output <= "11110101";
when "0010000100" => output <= "11110010";
when "0010000101" => output <= "11101111";
when "0010000110" => output <= "11101100";
when "0010000111" => output <= "11101001";
when "0010001000" => output <= "11100110";
when "0010001001" => output <= "11100011";
when "0010001010" => output <= "11100000";
when "0010001011" => output <= "11011101";
when "0010001100" => output <= "11011010";
when "0010001101" => output <= "11010111";
when "0010001110" => output <= "11010100";
when "0010001111" => output <= "11010001";
when "0010010000" => output <= "11001110";
when "0010010001" => output <= "11001011";
when "0010010010" => output <= "11001000";
when "0010010011" => output <= "11000101";
when "0010010100" => output <= "11000011";
when "0010010101" => output <= "11000000";
when "0010010110" => output <= "10111101";
when "0010010111" => output <= "10111010";
when "0010011000" => output <= "10111000";
when "0010011001" => output <= "10110101";
when "0010011010" => output <= "10110011";
when "0010011011" => output <= "10110000";
when "0010011100" => output <= "10101110";
when "0010011101" => output <= "10101011";
when "0010011110" => output <= "10101001";
when "0010011111" => output <= "10100111";
when "0010100000" => output <= "10100101";
when "0010100001" => output <= "10100010";
when "0010100010" => output <= "10100000";
when "0010100011" => output <= "10011110";
when "0010100100" => output <= "10011100";
when "0010100101" => output <= "10011010";
when "0010100110" => output <= "10011000";
when "0010100111" => output <= "10010111";
when "0010101000" => output <= "10010101";
when "0010101001" => output <= "10010011";
when "0010101010" => output <= "10010010";
when "0010101011" => output <= "10010000";
when "0010101100" => output <= "10001111";
when "0010101101" => output <= "10001101";
when "0010101110" => output <= "10001100";
when "0010101111" => output <= "10001011";
when "0010110000" => output <= "10001001";
when "0010110001" => output <= "10001000";
when "0010110010" => output <= "10000111";
when "0010110011" => output <= "10000110";
when "0010110100" => output <= "10000101";
when "0010110101" => output <= "10000101";
when "0010110110" => output <= "10000100";
when "0010110111" => output <= "10000011";
when "0010111000" => output <= "10000011";
when "0010111001" => output <= "10000010";
when "0010111010" => output <= "10000010";
when "0010111011" => output <= "10000001";
when "0010111100" => output <= "10000001";
when "0010111101" => output <= "10000001";
when "0010111110" => output <= "10000001";
when "0010111111" => output <= "10000001";
when "0011000000" => output <= "10000001";
when "0011000001" => output <= "10000001";
when "0011000010" => output <= "10000001";
when "0011000011" => output <= "10000001";
when "0011000100" => output <= "10000001";
when "0011000101" => output <= "10000010";
when "0011000110" => output <= "10000010";
when "0011000111" => output <= "10000011";
when "0011001000" => output <= "10000011";
when "0011001001" => output <= "10000100";
when "0011001010" => output <= "10000101";
when "0011001011" => output <= "10000110";
when "0011001100" => output <= "10000111";
when "0011001101" => output <= "10001000";
when "0011001110" => output <= "10001001";
when "0011001111" => output <= "10001010";
when "0011010000" => output <= "10001011";
when "0011010001" => output <= "10001101";
when "0011010010" => output <= "10001110";
when "0011010011" => output <= "10001111";
when "0011010100" => output <= "10010001";
when "0011010101" => output <= "10010010";
when "0011010110" => output <= "10010100";
when "0011010111" => output <= "10010110";
when "0011011000" => output <= "10011000";
when "0011011001" => output <= "10011001";
when "0011011010" => output <= "10011011";
when "0011011011" => output <= "10011101";
when "0011011100" => output <= "10011111";
when "0011011101" => output <= "10100001";
when "0011011110" => output <= "10100100";
when "0011011111" => output <= "10100110";
when "0011100000" => output <= "10101000";
when "0011100001" => output <= "10101010";
when "0011100010" => output <= "10101101";
when "0011100011" => output <= "10101111";
when "0011100100" => output <= "10110001";
when "0011100101" => output <= "10110100";
when "0011100110" => output <= "10110111";
when "0011100111" => output <= "10111001";
when "0011101000" => output <= "10111100";
when "0011101001" => output <= "10111110";
when "0011101010" => output <= "11000001";
when "0011101011" => output <= "11000100";
when "0011101100" => output <= "11000111";
when "0011101101" => output <= "11001010";
when "0011101110" => output <= "11001100";
when "0011101111" => output <= "11001111";
when "0011110000" => output <= "11010010";
when "0011110001" => output <= "11010101";
when "0011110010" => output <= "11011000";
when "0011110011" => output <= "11011011";
when "0011110100" => output <= "11011110";
when "0011110101" => output <= "11100001";
when "0011110110" => output <= "11100100";
when "0011110111" => output <= "11100111";
when "0011111000" => output <= "11101011";
when "0011111001" => output <= "11101110";
when "0011111010" => output <= "11110001";
when "0011111011" => output <= "11110100";
when "0011111100" => output <= "11110111";
when "0011111101" => output <= "11111010";
when "0011111110" => output <= "11111101";

-- triangle wave
when "0100000000" => output <= "00000000";
when "0100000001" => output <= "00000010";
when "0100000010" => output <= "00000100";
when "0100000011" => output <= "00000110";
when "0100000100" => output <= "00001000";
when "0100000101" => output <= "00001010";
when "0100000110" => output <= "00001100";
when "0100000111" => output <= "00001110";
when "0100001000" => output <= "00010000";
when "0100001001" => output <= "00010010";
when "0100001010" => output <= "00010100";
when "0100001011" => output <= "00010110";
when "0100001100" => output <= "00011000";
when "0100001101" => output <= "00011010";
when "0100001110" => output <= "00011100";
when "0100001111" => output <= "00011110";
when "0100010000" => output <= "00100000";
when "0100010001" => output <= "00100010";
when "0100010010" => output <= "00100100";
when "0100010011" => output <= "00100110";
when "0100010100" => output <= "00101000";
when "0100010101" => output <= "00101010";
when "0100010110" => output <= "00101100";
when "0100010111" => output <= "00101110";
when "0100011000" => output <= "00110000";
when "0100011001" => output <= "00110010";
when "0100011010" => output <= "00110100";
when "0100011011" => output <= "00110110";
when "0100011100" => output <= "00111000";
when "0100011101" => output <= "00111010";
when "0100011110" => output <= "00111100";
when "0100011111" => output <= "00111110";
when "0100100000" => output <= "01000000";
when "0100100001" => output <= "01000010";
when "0100100010" => output <= "01000100";
when "0100100011" => output <= "01000110";
when "0100100100" => output <= "01001000";
when "0100100101" => output <= "01001010";
when "0100100110" => output <= "01001100";
when "0100100111" => output <= "01001110";
when "0100101000" => output <= "01010000";
when "0100101001" => output <= "01010010";
when "0100101010" => output <= "01010100";
when "0100101011" => output <= "01010110";
when "0100101100" => output <= "01011000";
when "0100101101" => output <= "01011010";
when "0100101110" => output <= "01011100";
when "0100101111" => output <= "01011110";
when "0100110000" => output <= "01100000";
when "0100110001" => output <= "01100010";
when "0100110010" => output <= "01100100";
when "0100110011" => output <= "01100110";
when "0100110100" => output <= "01101000";
when "0100110101" => output <= "01101010";
when "0100110110" => output <= "01101100";
when "0100110111" => output <= "01101110";
when "0100111000" => output <= "01110000";
when "0100111001" => output <= "01110010";
when "0100111010" => output <= "01110100";
when "0100111011" => output <= "01110110";
when "0100111100" => output <= "01111000";
when "0100111101" => output <= "01111010";
when "0100111110" => output <= "01111100";
when "0100111111" => output <= "01111110";
when "0101000000" => output <= "01111111";
when "0101000001" => output <= "01111101";
when "0101000010" => output <= "01111011";
when "0101000011" => output <= "01111001";
when "0101000100" => output <= "01110111";
when "0101000101" => output <= "01110101";
when "0101000110" => output <= "01110011";
when "0101000111" => output <= "01110001";
when "0101001000" => output <= "01101111";
when "0101001001" => output <= "01101101";
when "0101001010" => output <= "01101011";
when "0101001011" => output <= "01101001";
when "0101001100" => output <= "01100111";
when "0101001101" => output <= "01100101";
when "0101001110" => output <= "01100011";
when "0101001111" => output <= "01100001";
when "0101010000" => output <= "01011111";
when "0101010001" => output <= "01011101";
when "0101010010" => output <= "01011011";
when "0101010011" => output <= "01011001";
when "0101010100" => output <= "01010111";
when "0101010101" => output <= "01010101";
when "0101010110" => output <= "01010011";
when "0101010111" => output <= "01010001";
when "0101011000" => output <= "01001111";
when "0101011001" => output <= "01001101";
when "0101011010" => output <= "01001011";
when "0101011011" => output <= "01001001";
when "0101011100" => output <= "01000111";
when "0101011101" => output <= "01000101";
when "0101011110" => output <= "01000011";
when "0101011111" => output <= "01000001";
when "0101100000" => output <= "00111111";
when "0101100001" => output <= "00111101";
when "0101100010" => output <= "00111011";
when "0101100011" => output <= "00111001";
when "0101100100" => output <= "00110111";
when "0101100101" => output <= "00110101";
when "0101100110" => output <= "00110011";
when "0101100111" => output <= "00110001";
when "0101101000" => output <= "00101111";
when "0101101001" => output <= "00101101";
when "0101101010" => output <= "00101011";
when "0101101011" => output <= "00101001";
when "0101101100" => output <= "00100111";
when "0101101101" => output <= "00100101";
when "0101101110" => output <= "00100011";
when "0101101111" => output <= "00100001";
when "0101110000" => output <= "00011111";
when "0101110001" => output <= "00011101";
when "0101110010" => output <= "00011011";
when "0101110011" => output <= "00011001";
when "0101110100" => output <= "00010111";
when "0101110101" => output <= "00010101";
when "0101110110" => output <= "00010011";
when "0101110111" => output <= "00010001";
when "0101111000" => output <= "00001111";
when "0101111001" => output <= "00001101";
when "0101111010" => output <= "00001011";
when "0101111011" => output <= "00001001";
when "0101111100" => output <= "00000111";
when "0101111101" => output <= "00000101";
when "0101111110" => output <= "00000011";
when "0101111111" => output <= "00000001";
when "0110000000" => output <= "11111111";
when "0110000001" => output <= "11111101";
when "0110000010" => output <= "11111011";
when "0110000011" => output <= "11111001";
when "0110000100" => output <= "11110111";
when "0110000101" => output <= "11110101";
when "0110000110" => output <= "11110011";
when "0110000111" => output <= "11110001";
when "0110001000" => output <= "11101111";
when "0110001001" => output <= "11101101";
when "0110001010" => output <= "11101011";
when "0110001011" => output <= "11101001";
when "0110001100" => output <= "11100111";
when "0110001101" => output <= "11100101";
when "0110001110" => output <= "11100011";
when "0110001111" => output <= "11100001";
when "0110010000" => output <= "11011111";
when "0110010001" => output <= "11011101";
when "0110010010" => output <= "11011011";
when "0110010011" => output <= "11011001";
when "0110010100" => output <= "11010111";
when "0110010101" => output <= "11010101";
when "0110010110" => output <= "11010011";
when "0110010111" => output <= "11010001";
when "0110011000" => output <= "11001111";
when "0110011001" => output <= "11001101";
when "0110011010" => output <= "11001011";
when "0110011011" => output <= "11001001";
when "0110011100" => output <= "11000111";
when "0110011101" => output <= "11000101";
when "0110011110" => output <= "11000011";
when "0110011111" => output <= "11000001";
when "0110100000" => output <= "10111111";
when "0110100001" => output <= "10111101";
when "0110100010" => output <= "10111011";
when "0110100011" => output <= "10111001";
when "0110100100" => output <= "10110111";
when "0110100101" => output <= "10110101";
when "0110100110" => output <= "10110011";
when "0110100111" => output <= "10110001";
when "0110101000" => output <= "10101111";
when "0110101001" => output <= "10101101";
when "0110101010" => output <= "10101011";
when "0110101011" => output <= "10101001";
when "0110101100" => output <= "10100111";
when "0110101101" => output <= "10100101";
when "0110101110" => output <= "10100011";
when "0110101111" => output <= "10100001";
when "0110110000" => output <= "10011111";
when "0110110001" => output <= "10011101";
when "0110110010" => output <= "10011011";
when "0110110011" => output <= "10011001";
when "0110110100" => output <= "10010111";
when "0110110101" => output <= "10010101";
when "0110110110" => output <= "10010011";
when "0110110111" => output <= "10010001";
when "0110111000" => output <= "10001111";
when "0110111001" => output <= "10001101";
when "0110111010" => output <= "10001011";
when "0110111011" => output <= "10001001";
when "0110111100" => output <= "10000111";
when "0110111101" => output <= "10000101";
when "0110111110" => output <= "10000011";
when "0110111111" => output <= "10000001";
when "0111000000" => output <= "10000010";
when "0111000001" => output <= "10000100";
when "0111000010" => output <= "10000110";
when "0111000011" => output <= "10001000";
when "0111000100" => output <= "10001010";
when "0111000101" => output <= "10001100";
when "0111000110" => output <= "10001110";
when "0111000111" => output <= "10010000";
when "0111001000" => output <= "10010010";
when "0111001001" => output <= "10010100";
when "0111001010" => output <= "10010110";
when "0111001011" => output <= "10011000";
when "0111001100" => output <= "10011010";
when "0111001101" => output <= "10011100";
when "0111001110" => output <= "10011110";
when "0111001111" => output <= "10100000";
when "0111010000" => output <= "10100010";
when "0111010001" => output <= "10100100";
when "0111010010" => output <= "10100110";
when "0111010011" => output <= "10101000";
when "0111010100" => output <= "10101010";
when "0111010101" => output <= "10101100";
when "0111010110" => output <= "10101110";
when "0111010111" => output <= "10110000";
when "0111011000" => output <= "10110010";
when "0111011001" => output <= "10110100";
when "0111011010" => output <= "10110110";
when "0111011011" => output <= "10111000";
when "0111011100" => output <= "10111010";
when "0111011101" => output <= "10111100";
when "0111011110" => output <= "10111110";
when "0111011111" => output <= "11000000";
when "0111100000" => output <= "11000010";
when "0111100001" => output <= "11000100";
when "0111100010" => output <= "11000110";
when "0111100011" => output <= "11001000";
when "0111100100" => output <= "11001010";
when "0111100101" => output <= "11001100";
when "0111100110" => output <= "11001110";
when "0111100111" => output <= "11010000";
when "0111101000" => output <= "11010010";
when "0111101001" => output <= "11010100";
when "0111101010" => output <= "11010110";
when "0111101011" => output <= "11011000";
when "0111101100" => output <= "11011010";
when "0111101101" => output <= "11011100";
when "0111101110" => output <= "11011110";
when "0111101111" => output <= "11100000";
when "0111110000" => output <= "11100010";
when "0111110001" => output <= "11100100";
when "0111110010" => output <= "11100110";
when "0111110011" => output <= "11101000";
when "0111110100" => output <= "11101010";
when "0111110101" => output <= "11101100";
when "0111110110" => output <= "11101110";
when "0111110111" => output <= "11110000";
when "0111111000" => output <= "11110010";
when "0111111001" => output <= "11110100";
when "0111111010" => output <= "11110110";
when "0111111011" => output <= "11111000";
when "0111111100" => output <= "11111010";
when "0111111101" => output <= "11111100";
when "0111111110" => output <= "11111110";

when others => output <= (others => '0');
end case;

end process;

end;